// Bradyn Hinman
// 3/15/2023
// Skeeball Display

module skeeballDisplay(state, score, HEX5, HEX4, HEX3, HEX2, HEX1, HEX0);
	input [1:0] state;
	input [6:0] score;
	output [6:0] HEX5, HEX4, HEX3, HEX2, HEX1, HEX0;
	
	
	
	
endmodule