// Bradyn Hinman
// 3/15/2023
// Skeeball State Machine

module skeeballState(state, balls, display);
	output [1:0] state;
	output [8:0] balls;
	output [41:0] display;
	
	reg [6:0] gamescore, highscore;
	
	
endmodule